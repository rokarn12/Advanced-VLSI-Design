parameter int NUM_TAPS = 170;
parameter logic signed [15:0] fir_coefs[0:NUM_TAPS-1] = '{
    16'b0000000000000000,
    16'b1111111111111000,
    16'b1111111111101010,
    16'b1111111111010010,
    16'b1111111110101111,
    16'b1111111110000101,
    16'b1111111101011100,
    16'b1111111100111101,
    16'b1111111100110100,
    16'b1111111101000110,
    16'b1111111101110101,
    16'b1111111110111010,
    16'b0000000000000110,
    16'b0000000001000111,
    16'b0000000001101100,
    16'b0000000001101011,
    16'b0000000001000110,
    16'b0000000000001011,
    16'b1111111111001110,
    16'b1111111110100101,
    16'b1111111110100000,
    16'b1111111111000000,
    16'b1111111111111010,
    16'b0000000000110111,
    16'b0000000001100000,
    16'b0000000001100011,
    16'b0000000000111101,
    16'b1111111111111100,
    16'b1111111110111001,
    16'b1111111110010001,
    16'b1111111110010101,
    16'b1111111111000111,
    16'b0000000000010100,
    16'b0000000001011110,
    16'b0000000010000100,
    16'b0000000001110110,
    16'b0000000000110100,
    16'b1111111111010111,
    16'b1111111110000101,
    16'b1111111101100001,
    16'b1111111101111111,
    16'b1111111111010110,
    16'b0000000001000111,
    16'b0000000010100001,
    16'b0000000010111110,
    16'b0000000010001011,
    16'b0000000000011000,
    16'b1111111110010010,
    16'b1111111100110000,
    16'b1111111100011111,
    16'b1111111101101110,
    16'b0000000000000011,
    16'b0000000010100100,
    16'b0000000100001100,
    16'b0000000100001001,
    16'b0000000010010011,
    16'b1111111111010010,
    16'b1111111100010010,
    16'b1111111010101000,
    16'b1111111011001001,
    16'b1111111101110101,
    16'b0000000001110000,
    16'b0000000101010101,
    16'b0000000110111110,
    16'b0000000101101111,
    16'b0000000001110100,
    16'b1111111100101000,
    16'b1111111000010000,
    16'b1111110110101110,
    16'b1111111001001000,
    16'b1111111110111110,
    16'b0000000110001101,
    16'b0000001011111001,
    16'b0000001101001101,
    16'b0000001000101111,
    16'b1111111111010000,
    16'b1111110011110010,
    16'b1111101010111111,
    16'b1111101001100010,
    16'b1111110010101001,
    16'b0000000110101100,
    16'b0000100010101100,
    16'b0001000000111101,
    16'b0001011010100000,
    16'b0001101001000111,
    16'b0001101001000111,
    16'b0001011010100000,
    16'b0001000000111101,
    16'b0000100010101100,
    16'b0000000110101100,
    16'b1111110010101001,
    16'b1111101001100010,
    16'b1111101010111111,
    16'b1111110011110010,
    16'b1111111111010000,
    16'b0000001000101111,
    16'b0000001101001101,
    16'b0000001011111001,
    16'b0000000110001101,
    16'b1111111110111110,
    16'b1111111001001000,
    16'b1111110110101110,
    16'b1111111000010000,
    16'b1111111100101000,
    16'b0000000001110100,
    16'b0000000101101111,
    16'b0000000110111110,
    16'b0000000101010101,
    16'b0000000001110000,
    16'b1111111101110101,
    16'b1111111011001001,
    16'b1111111010101000,
    16'b1111111100010010,
    16'b1111111111010010,
    16'b0000000010010011,
    16'b0000000100001001,
    16'b0000000100001100,
    16'b0000000010100100,
    16'b0000000000000011,
    16'b1111111101101110,
    16'b1111111100011111,
    16'b1111111100110000,
    16'b1111111110010010,
    16'b0000000000011000,
    16'b0000000010001011,
    16'b0000000010111110,
    16'b0000000010100001,
    16'b0000000001000111,
    16'b1111111111010110,
    16'b1111111101111111,
    16'b1111111101100001,
    16'b1111111110000101,
    16'b1111111111010111,
    16'b0000000000110100,
    16'b0000000001110110,
    16'b0000000010000100,
    16'b0000000001011110,
    16'b0000000000010100,
    16'b1111111111000111,
    16'b1111111110010101,
    16'b1111111110010001,
    16'b1111111110111001,
    16'b1111111111111100,
    16'b0000000000111101,
    16'b0000000001100011,
    16'b0000000001100000,
    16'b0000000000110111,
    16'b1111111111111010,
    16'b1111111111000000,
    16'b1111111110100000,
    16'b1111111110100101,
    16'b1111111111001110,
    16'b0000000000001011,
    16'b0000000001000110,
    16'b0000000001101011,
    16'b0000000001101100,
    16'b0000000001000111,
    16'b0000000000000110,
    16'b1111111110111010,
    16'b1111111101110101,
    16'b1111111101000110,
    16'b1111111100110100,
    16'b1111111100111101,
    16'b1111111101011100,
    16'b1111111110000101,
    16'b1111111110101111,
    16'b1111111111010010,
    16'b1111111111101010,
    16'b1111111111111000,
    16'b0000000000000000
};
