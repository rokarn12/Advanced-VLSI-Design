// Definitions for scalability
`define VMEM_SPACE 64
`define VMEM_BITS 6

`define PMEM_SPACE 32
`define PMEM_BITS 5

`define VPN_WIDTH 6

`define PPN_WIDTH 4

`define OFFSET_WIDTH 2

`define NUM_PHYS_PAGES 8
